library ieee ;
    use ieee.std_logic_1164.all ;
    use ieee.numeric_std.all ;

entity compteur is
    port (
        clock, raz, en_count: in std_logic;
        
    ) ;
end compteur ; 

architecture arch_compteur of compteur is

begin

end architecture ;